//Modified from ARA SRAM
